`timescale 1ns / 1ps

module debouncher(
    input clk,
    input pbin,     
    output pbout  
    );

  

endmodule
