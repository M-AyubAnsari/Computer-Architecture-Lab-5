`timescale 1ns / 1ps
module debouncer(
    input clk,
    input pbin,
    output pbout
    );
endmodule
